class packet
  // write your code.
endclass: check
