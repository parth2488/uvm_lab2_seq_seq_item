
class packet_sequence.sv

  // Add your code here.
  // bhen da takas... 
  
endclass : checck

